--
-- VHDL Architecture my_project1_lib.Reg.Behavior
--
-- Created:
--          by - powel.UNKNOWN (LAPTOP-627UE0BV)
--          at - 13:12:02 01/28/2019
--
-- using Mentor Graphics HDL Designer(TM) 2015.1b (Build 4)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Reg IS
  GENERIC(width : NATURAL RANGE 1 to 64 := 8);
  PORT(D : IN std_ulogic_vector(width - 1 DOWNTO 0);
    Q : OUT std_ulogic_vector(width - 1 DOWNTO 0);
    clk, enable, rst : IN std_ulogic);
END ENTITY Reg;

--
ARCHITECTURE Behavior OF Reg IS
BEGIN
  PROCESS(D, clk, enable, rst)
    CONSTANT zero : std_ulogic_vector(width - 1 DOWNTO 0) := (others => '0');
    
  BEGIN
    IF(rising_edge(clk) AND enable = '1') THEN
      Q <= D;
    END IF;
    IF(rst = '1') THEN
      Q <= zero;
    END IF;
  END PROCESS;
END ARCHITECTURE Behavior;

